// 7-bit Mastrovito multiplier
// Primitive polynomial to use: x^7 + x + 1

module Mastrovito7(a, b, c);
endmodule