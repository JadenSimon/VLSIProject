module PointMultiplier(point, scalar, clk) 


endmodule 