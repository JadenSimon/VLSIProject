// 7-bit Mastrovito multiplier
// Primitive polynomial to use: x^7 + x + 1
// Resources: 
// https://pdfs.semanticscholar.org/501f/856a68c5231d93c82ce89456bff55842b13b.pdf
// https://online.tugraz.at/tug_online/voe_main2.getvolltext?pCurrPk=43036

module Mastrovito7(a, b, c);
endmodule